library verilog;
use verilog.vl_types.all;
entity lab_parteA_vlg_check_tst is
    port(
        LED             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab_parteA_vlg_check_tst;
