library verilog;
use verilog.vl_types.all;
entity ParteC_vlg_vec_tst is
end ParteC_vlg_vec_tst;
