library verilog;
use verilog.vl_types.all;
entity lab_parteA_vlg_vec_tst is
end lab_parteA_vlg_vec_tst;
